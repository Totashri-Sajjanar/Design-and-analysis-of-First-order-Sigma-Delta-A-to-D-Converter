* C:\Users\Lenovo\eSim-Workspace\Sigma_DeltaAdc\Sigma_DeltaAdc1.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 10/07/22 00:56:58

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U5  Comp_out Clk GND Dlatch_out d_latch		
v2  Analog_in GND pulse		
v4  Clk GND pulse		
SC1  Analog_in Net-_SC1-Pad2_ sky130_fd_pr__cap_mim_m3_1		
v3  Net-_X1-Pad1_ Net-_X1-Pad2_ DC		
X1  Net-_X1-Pad1_ Net-_X1-Pad2_ Net-_SC1-Pad2_ Net-_U4-Pad2_ Dif_out GND avsd_opamp		
SC2  Net-_SC1-Pad2_ Dif_out Net-_SC2-Pad3_ sky130_fd_pr__res_generic_pd		
SC3  Dif_out Net-_SC3-Pad2_ Net-_SC2-Pad3_ sky130_fd_pr__res_generic_pd		
X2  Net-_X2-Pad1_ Net-_X2-Pad2_ GND Net-_SC3-Pad2_ Intg_out GND avsd_opamp		
v5  Net-_X2-Pad1_ Net-_X2-Pad2_ DC		
X3  Net-_X3-Pad1_ Net-_X3-Pad2_ ? GND Comp_out GND avsd_opamp		
v6  Net-_X3-Pad1_ Net-_X3-Pad2_ DC		
U9  Dlatch_out Bit_out adc_bridge_1		
U4  Bit_out Net-_U4-Pad2_ dac_bridge_1		
v1  Net-_SC2-Pad3_ GND DC		
U1  Analog_in plot_v1		
U2  Clk plot_v1		
U3  Dif_out plot_v1		
U6  Intg_out plot_v1		
U7  Comp_out plot_v1		
U8  Dlatch_out plot_v1		
U10  Bit_out plot_v1		
SC4  Net-_SC3-Pad2_ Intg_out sky130_fd_pr__cap_mim_m3_1		
scmode1  SKY130mode		

.end
