* C:\Users\Lenovo\eSim-Workspace\Sigma_DeltaAdc\Sigma_DeltaAdc2.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 10/07/22 01:15:38

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U5  Comp_out Clk GND Dlatch_out d_latch		
v2  Analog_in GND pulse		
v4  Clk GND pulse		
v3  Net-_X1-Pad1_ Net-_X1-Pad2_ DC		
X1  Net-_X1-Pad1_ Net-_X1-Pad2_ Net-_C1-Pad2_ Net-_U4-Pad2_ Dif_out GND avsd_opamp		
X2  Net-_X2-Pad1_ Net-_X2-Pad2_ GND Net-_C2-Pad2_ Intg_out GND avsd_opamp		
v5  Net-_X2-Pad1_ Net-_X2-Pad2_ DC		
X3  Net-_X3-Pad1_ Net-_X3-Pad2_ ? GND Comp_out GND avsd_opamp		
v6  Net-_X3-Pad1_ Net-_X3-Pad2_ DC		
U9  Dlatch_out Bit_out adc_bridge_1		
U4  Bit_out Net-_U4-Pad2_ dac_bridge_1		
U1  Analog_in plot_v1		
U2  Clk plot_v1		
U3  Dif_out plot_v1		
U6  Intg_out plot_v1		
U7  Comp_out plot_v1		
U8  Dlatch_out plot_v1		
U10  Bit_out plot_v1		
scmode1  SKY130mode		
R1  Net-_C1-Pad2_ Dif_out 1000		
R2  Dif_out Net-_C2-Pad2_ 1000		
C1  Analog_in Net-_C1-Pad2_ 1p		
C2  Intg_out Net-_C2-Pad2_ 1p		

.end
